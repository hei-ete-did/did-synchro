PACKAGE Common IS

  function requiredBitNb (val : integer) return integer;

END Common;
